`include "3_VideoSync_Generator.v"

module test_hvsync_top(clk, reset, hsync, vsync, rgb);

  input clk, reset;
  output hsync, vsync;
  output [2:0] rgb;
  
  wire display_on;
  wire [8:0] hpos;
  wire [8:0] vpos;

  hvsync_generator hvsync_gen(
    .clk(clk),
    .reset(0),
    .hsync(hsync),
    .vsync(vsync),
    .display_on(display_on),
    .hpos(hpos),
    .vpos(vpos)
  );

  wire r = display_on & (((hpos&7)==0) | ((vpos&7)==0));
  wire g = display_on & vpos[4];
  wire b = display_on & hpos[4];

  assign rgb = {b, g, r};

endmodule
